`default_nettype none
`include "clockworks.v"
`include "emitter_uart.v"

module Memory (
    input              clk,
    input      [31:0]  mem_addr,  // address to be read
    output reg [31:0]  mem_rdata, // data read from memory
    input   	         mem_rstrb,  // goes high when processor wants to read
    input      [31:0]  mem_wdata,
    input      [3:0]   mem_wmask
);

  reg [31:0] MEM [0:1535]; 

`ifdef BENCH
  localparam slow_bit=12;
`else
  localparam slow_bit=17;
`endif

  // Memory-mapped IO in IO page, 1-hot addressing in word address.   
  localparam IO_LEDS_bit      = 0;  // W five leds - offset = 32'h400004
  localparam IO_UART_DAT_bit  = 1;  // W data to send (8 bits), offset = 32'h400008
  localparam IO_UART_CNTL_bit = 2;  // R status. bit 9: busy sending, offset = 32'h400010

  // Converts an IO_xxx_bit constant into an offset in IO page.
  function [31:0] IO_BIT_TO_OFFSET;
    input [31:0] bitid;
    begin
      IO_BIT_TO_OFFSET = 1 << (bitid + 2);
    end
  endfunction

`include "riscv_assembly.v"
   integer    L0_      = 12;
   integer    L1_      = 20;
   integer    L2_      = 52;      
   integer    wait_    = 104;
   integer    wait_L0_ = 112;
   integer    putc_    = 124; 
   integer    putc_L0_ = 132;
   
   initial begin
      LI(sp,32'h1800);   // End of RAM, 6kB
      LI(gp,32'h400000); // IO page

   Label(L0_);

      // Count from 0 to 15 on the LEDs      
      LI(s0,16); // upper bound of loop
      LI(a0,0);
   Label(L1_);
      SW(a0,gp,IO_BIT_TO_OFFSET(IO_LEDS_bit));
      CALL(LabelRef(wait_));
      ADDI(a0,a0,1);
      BNE(a0,s0,LabelRef(L1_));

      // Send abcdef...xyz to the UART
      LI(s0,26); // upper bound of loop     
      LI(a0,"a");
      LI(s1,0);
   Label(L2_);
      CALL(LabelRef(putc_));
      ADDI(a0,a0,1);
      ADDI(s1,s1,1);
      BNE(s1,s0,LabelRef(L2_));

      // CR;LF
      LI(a0,13);
      CALL(LabelRef(putc_));
      LI(a0,10);
      CALL(LabelRef(putc_));
      
      J(LabelRef(L0_));
      
      EBREAK(); // I systematically keep it before functions
                // in case I decide to remove the loop...

   Label(wait_);
      LI(t0,1);
      SLLI(t0,t0,slow_bit);
   Label(wait_L0_);
      ADDI(t0,t0,-1);
      BNEZ(t0,LabelRef(wait_L0_));
      RET();

   Label(putc_);
      // Send character to UART
      SW(a0,gp,IO_BIT_TO_OFFSET(IO_UART_DAT_bit));
      // Read UART status, and loop until bit 9 (busy sending)
      // is zero.
      LI(t0,1<<9);
   Label(putc_L0_);
      LW(t1,gp,IO_BIT_TO_OFFSET(IO_UART_CNTL_bit));     
      AND(t1,t1,t0);
      BNEZ(t1,LabelRef(putc_L0_));
      RET();
	   
      endASM();
   end

  wire [29:0] word_addr = mem_addr[31:2];
  always @(posedge clk) begin
    if(mem_rstrb) begin
      mem_rdata <= MEM[mem_addr[31:2]];
    end
    if (mem_wmask[0]) MEM[word_addr][7:0  ] <= mem_wdata[7:0  ];
    if (mem_wmask[1]) MEM[word_addr][15:8 ] <= mem_wdata[15:8 ];
    if (mem_wmask[2]) MEM[word_addr][23:16] <= mem_wdata[23:16];
    if (mem_wmask[3]) MEM[word_addr][31:24] <= mem_wdata[31:24];
  end
endmodule

module Processor (
    input 	          clk,
    input 	          resetn,
    output     [31:0] mem_addr, 
    input      [31:0] mem_rdata, 
    output 	          mem_rstrb,
    output     [31:0] mem_wdata,
    output     [3:0]  mem_wmask
);

  reg [31:0] PC=0;
  reg [31:0] instr;

  // decoder
  // R-type  [31  funct7     25]  [24  rs2  20]  [19  rs1  15]  [14  funct3  12]  [11  rd        7]  [6  opcode  0]
  // S-type  [31  imm[11:5]  25]  [24  rs2  20]  [19  rs1  15]  [14  funct3  12]  [11  imm[4:0]  7]  [6  opcode  0]
  // I-type  [31  imm[11:0]                 20]  [19  rs1  15]  [14  funct3  12]  [11  rd        7]  [6  opcode  0]
  // U-type  [31  imm[31:12]                                                 12]  [11  rd        7]  [6  opcode  0]

  // decode op codes
  wire isALUreg  =  (instr[6:0] == 7'b0110011); // rd <- rs1 OP rs2   
  wire isALUimm  =  (instr[6:0] == 7'b0010011); // rd <- rs1 OP Iimm
  wire isBranch  =  (instr[6:0] == 7'b1100011); // if(rs1 OP rs2) PC<-PC+Bimm
  wire isJALR    =  (instr[6:0] == 7'b1100111); // rd <- PC+4; PC<-rs1+Iimm
  wire isJAL     =  (instr[6:0] == 7'b1101111); // rd <- PC+4; PC<-PC+Jimm
  wire isAUIPC   =  (instr[6:0] == 7'b0010111); // rd <- PC + Uimm
  wire isLUI     =  (instr[6:0] == 7'b0110111); // rd <- Uimm   
  wire isLoad    =  (instr[6:0] == 7'b0000011); // rd <- mem[rs1+Iimm]
  wire isStore   =  (instr[6:0] == 7'b0100011); // mem[rs1+Simm] <- rs2
  wire isSYSTEM  =  (instr[6:0] == 7'b1110011); // special

  // decode source and destination registers
  wire [4:0] rs2Id = instr[24:20];
  wire [4:0] rs1Id = instr[19:15];
  wire [4:0] rdId  = instr[11:7];

  // extract funct7 and funct3
  wire [6:0] funct7 = instr[31:25];
  wire [2:0] funct3 = instr[14:12];

  // build immediates for each instruction type
  wire [31:0] Uimm={    instr[31],   instr[30:12], {12{1'b0}}};
  wire [31:0] Iimm={{21{instr[31]}}, instr[30:20]};
  wire [31:0] Simm={{21{instr[31]}}, instr[30:25], instr[11:7]};
  wire [31:0] Bimm={{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0};
  wire [31:0] Jimm={{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};

  // register bank
  reg [31:0] RegisterBank [0:31];
  reg [31:0] rs1;
  reg [31:0] rs2;
  wire [31:0] writeBackData;
  wire writeBackEn;

  `ifdef BENCH   
    integer     i;
    initial begin
      for(i=0; i<32; ++i) begin
        RegisterBank[i] = 0;
      end
    end
  `endif   

  // ALU
  wire [31:0] aluIn1 = rs1;
  wire [31:0] aluIn2 = isALUreg | isBranch ? rs2 : Iimm;
  reg [31:0] aluOut;
  wire [4:0] shamt = isALUreg ? rs2[4:0] : instr[24:20]; // shift amount

  wire [31:0] aluPlus = aluIn1 + aluIn2;
  wire [32:0] aluMinus = {1'b1, ~aluIn2} + {1'b0, aluIn1} + 33'b1; // A-B = A + ~B + 1
  wire EQ = (aluMinus[31:0] == 0); // A==B if A-B = 0
  wire LTU = aluMinus[32]; // because aluMinus is sign extended, MSB 1 for negative
  wire LT = (aluIn1[31] ^ aluIn2[31]) ? aluIn1[31] : aluMinus[32]; // if signs differ then A < B if A is negative, else check if A-B is negative

  // Flip a 32 bit word. Used by the shifter (a single shifter for
  // left and right shifts, saves silicium !)
  function [31:0] flip32;
    input [31:0] x;
    flip32 = {x[ 0], x[ 1], x[ 2], x[ 3], x[ 4], x[ 5], x[ 6], x[ 7], 
		x[ 8], x[ 9], x[10], x[11], x[12], x[13], x[14], x[15], 
		x[16], x[17], x[18], x[19], x[20], x[21], x[22], x[23],
		x[24], x[25], x[26], x[27], x[28], x[29], x[30], x[31]};
  endfunction

  wire [31:0] shifter = $signed({instr[30] & aluIn1[31], shifter_in}) >>> aluIn2[4:0];
  wire [31:0] shifter_in = (funct3 == 3'b001) ? flip32(aluIn1) : aluIn1;
  wire [31:0] leftshift = flip32(shifter);

  // ADD/SUB/ADDI: funct7[5] 0=ADD, 1=SUB, instr[5]=I
  // SRL/SRLI/SRA/SRAI: funct7[5] 0=logical, 1=arthimetic
  always @(*) begin
    case (funct3)
      3'b000: aluOut = (funct7[5] & instr[5]) ? aluMinus[31:0] : aluPlus; // ADD/ADDI/SUB/SUBI
      3'b001: aluOut = leftshift;                                         // SLL
      3'b010: aluOut = {31'b0, LT};                                       // SLT
      3'b011: aluOut = {31'b0, LTU};                                      // SLTU
      3'b100: aluOut = (aluIn1 ^ aluIn2);                                 // XOR
      3'b101: aluOut = shifter;                                           // SRA/SRAI
      3'b110: aluOut = (aluIn1 | aluIn2);                                 // OR
      3'b111: aluOut = (aluIn1 & aluIn2);                                 // AND
    endcase
  end

  // The predicate for branch instructions
  reg takeBranch;
  always @(*) begin
    case(funct3)
      3'b000: takeBranch = EQ;
      3'b001: takeBranch = !EQ;
      3'b100: takeBranch = LT;
      3'b101: takeBranch = !LT;
      3'b110: takeBranch = LTU;
      3'b111: takeBranch = !LTU;
      default: takeBranch = 1'b0;
    endcase
  end

  wire [31:0] PCplusImm = PC + (instr[3] ? Jimm[31:0] :
                                instr[4] ? Uimm[31:0] :
                                Bimm);
  wire [31:0] PCplus4 = PC + 4;
  wire [31:0] nextPC = ((isBranch && takeBranch) || isJAL) ? PCplusImm :
                        isJALR ? {aluPlus[31:1], 1'b0} :
                        PCplus4;

  wire [31:0] loadstore_addr = rs1 + (isStore ? Simm : Iimm);

  // what will be written back to register
  assign writeBackData = (isJAL || isJALR)  ? PCplus4 :
                         isLUI              ? Uimm :
                         isAUIPC            ? PCplusImm :
                         isLoad             ? LOAD_data :
                                              aluOut;

  // are we writing back to a register (or somewhere else)
  assign writeBackEn = (state==EXECUTE && !isBranch && !isStore && !isLoad) || (state == WAIT_DATA); // save writeBackData to RegisterFile[rdId]


  // LOAD from memory                       
  wire mem_byteAccess = funct3[1:0] == 2'b00;
  wire mem_halfwordAccess = funct3[1:0] == 2'b01;

  wire [15:0] LOAD_halfword = loadstore_addr[1] ? mem_rdata[31:16] : mem_rdata[15:0];
  wire [15:0] LOAD_byte = loadstore_addr[0] ? LOAD_halfword[15:8] : LOAD_halfword[7:0];
  wire        LOAD_sign = !funct3[2] & (mem_byteAccess ? LOAD_byte[7] : LOAD_halfword[15]); // sign is MSB, or 0 if unsigned load (funct3==0)
  wire [31:0] LOAD_data = mem_byteAccess ? {{24{LOAD_sign}}, LOAD_byte} : mem_halfwordAccess ? {{16{LOAD_sign}}, LOAD_halfword} : mem_rdata;

  // STORE to memory
  assign mem_wdata[ 7: 0] = rs2[7:0];
  assign mem_wdata[15: 8] = loadstore_addr[0] ? rs2[7:0] : rs2[15: 8];
  assign mem_wdata[23:16] = loadstore_addr[1] ? rs2[7:0] : rs2[23:16];
  assign mem_wdata[31:24] = loadstore_addr[0] ? rs2[7:0] : loadstore_addr[1] ? rs2[15:8] : rs2[31:24];
  wire [3:0] STORE_wmask =
	      mem_byteAccess      ?
	            (loadstore_addr[1] ?
		          (loadstore_addr[0] ? 4'b1000 : 4'b0100) :
		          (loadstore_addr[0] ? 4'b0010 : 4'b0001)) :
	      mem_halfwordAccess ?
	            (loadstore_addr[1] ? 4'b1100 : 4'b0011) :
              4'b1111;

  // states
  // The state machine
  localparam FETCH_INSTR = 0;
  localparam WAIT_INSTR  = 1;
  localparam FETCH_REGS  = 2;
  localparam EXECUTE     = 3;
  localparam LOAD        = 4;
  localparam WAIT_DATA   = 5;
  localparam STORE       = 6;
  reg [2:0] state = FETCH_INSTR;

  // cycle
  always @(posedge clk) begin
    if (!resetn) begin
      PC <= 0;
      state <= FETCH_INSTR;
    end else begin
      if (writeBackEn && rdId != 0) begin
        RegisterBank[rdId] <= writeBackData;
        `ifdef BENCH	 
	        // $display("x%0d <= %b", rdId, writeBackData);
        `endif
      end;

      case (state)
        FETCH_INSTR: begin
          state <= WAIT_INSTR;
        end
        WAIT_INSTR: begin
          instr <= mem_rdata;
          state <= FETCH_REGS;
        end
        FETCH_REGS: begin
          rs1 <= RegisterBank[rs1Id];
          rs2 <= RegisterBank[rs2Id];
          state <= EXECUTE;
        end
        EXECUTE: begin
          if (!isSYSTEM) begin
            PC <= nextPC;
          end
          state <= isLoad ? LOAD : isStore ? STORE : FETCH_INSTR;
          `ifdef BENCH
            if(isSYSTEM) $finish();
          `endif
        end
        LOAD: begin
          state <= WAIT_DATA;
        end
        WAIT_DATA: begin
          state <= FETCH_INSTR;
        end
        STORE: begin
          state <= FETCH_INSTR;
        end
      endcase 
    end
  end

  // outputs
  assign mem_addr = (state == WAIT_INSTR || state == FETCH_INSTR) ? PC : loadstore_addr;
  assign mem_rstrb = (state == FETCH_INSTR || state == LOAD);
  assign mem_wmask = {4{(state == STORE)}} & STORE_wmask;

  `ifdef BENCH2
    always @(posedge clk) begin
      if (state == FETCH_REGS) begin
        case (1'b1)
          isALUreg: $display("ALUreg rd=%d rs1=%d rs2=%d funct3=%b", rdId, rs1Id, rs2Id, funct3);
          isALUimm: $display("ALUimm rd=%d rs1=%d imm=%0d funct3=%b", rdId, rs1Id, Iimm, funct3);
          isBranch: $display("BRANCH");
          isJAL:    $display("JAL");
          isJALR:   $display("JALR");
          isAUIPC:  $display("AUIPC");
          isLUI:    $display("LUI");	
          isLoad:   $display("LOAD");
          isStore:  $display("STORE");
          isSYSTEM: $display("SYSTEM");
        endcase
        if (isSYSTEM) $finish();
      end
    end
  `endif

endmodule

module SOC (
  input CLK,
  input RESET,
  output reg [4:0] LEDS,
  input RXD,
  output TXD
);

  wire clk;
  wire resetn;

  wire [31:0] mem_addr;
  wire [31:0] mem_rdata;
  wire mem_rstrb;
  wire [31:0] mem_wdata;
  wire [3:0]  mem_wmask;

//  Memory            |                   | Processor     
//                    |                   |                
//                    |  <<<<<<<<<<<<<<   | mem_addr                
//                    |  <<<<<<<<<<<<<<   | mem_rstrb                
//                    |  <<<<<<<<<<<<<<   | mem_wdata                
//                    |  <<<<<<<<<<<<<<   | mem_wmask   
//                    |                   |           
//          mem_rdata |  >> RAM_rdata >>  |                 
//                    |  >> IO_rdata  >>  |                 


  Processor CPU(
    .clk(clk),
    .resetn(resetn),
    .mem_rdata(mem_rdata), //input
    .mem_addr(mem_addr),   //output
    .mem_rstrb(mem_rstrb), //output
    .mem_wdata(mem_wdata), //output
    .mem_wmask(mem_wmask)  //output
  );

  wire [31:0] RAM_rdata;
  wire [29:0] mem_wordaddr = mem_addr[31:2];
  wire isIO  = mem_addr[22]; // 00000000000000000000000000000000
  wire isRAM = !isIO;
  wire mem_wstrb = |mem_wmask;

  Memory RAM(
    .clk(clk),
    .mem_addr(mem_addr),              //input
    .mem_rstrb(isRAM & mem_rstrb),    //input
    .mem_wdata(mem_wdata),            //input
    .mem_wmask({4{isRAM}}&mem_wmask), //input - if isIO will be 0000 to stop write to physical ram as addr is virtual only
    .mem_rdata(RAM_rdata)             //output
  );

  // virtual addresses
  // 00000000010000000000000000000000 = 0x400000  
  // 00000000010000000000000000000100 = 0x400004 = IO_LEDS_bit = 0
  // 00000000010000000000000000001000 = 0x400008 = IO_UART_DAT_BIT = 1
  // 00000000010000000000000000010000 = 0x400010 = IO_UART_CNTL_BIT = 2

  // mem_wordaddr = mem_addr[31:2];
  // 000000000100000000000000000001 = mem_wordaddr[IO_LEDS_bit] = 1
  // 000000000100000000000000000010 = mem_wordaddr[IO_UART_DAT_BIT] = 1
  // 000000000100000000000000000100 = mem_wordaddr[IO_UART_CNTL_BIT] = 1

  // Memory-mapped IO in IO page, 1-hot addressing in word address.   
  localparam IO_LEDS_bit      = 0;  // W five leds
  localparam IO_UART_DAT_bit  = 1;  // W data to send (8 bits) 
  localparam IO_UART_CNTL_bit = 2;  // R status. bit 9: busy sending
   
  always @(posedge clk) begin
    if(isIO & mem_wstrb & mem_wordaddr[IO_LEDS_bit]) begin
      LEDS <= mem_wdata;
    end
  end

  wire uart_valid = isIO & mem_wstrb & mem_wordaddr[IO_UART_DAT_bit];
  wire uart_ready;

  corescore_emitter_uart #(
    .clk_freq_hz(`CPU_FREQ*1000000),
    .baud_rate(1000000)			    
  ) UART(
    .i_clk(clk),
    .i_rst(!resetn),
    .i_data(mem_wdata[7:0]),
    .i_valid(uart_valid),
    .o_ready(uart_ready),
    .o_uart_tx(TXD)      			       
  );

     wire [31:0] IO_rdata = 
	       mem_wordaddr[IO_UART_CNTL_bit] ? { 22'b0, !uart_ready, 9'b0}
	                                      : 32'b0;
   
   assign mem_rdata = isRAM ? RAM_rdata : IO_rdata;

`ifdef BENCH
   always @(posedge clk) begin
      if(uart_valid) begin
	 $write("%c", mem_wdata[7:0] );
	 $fflush(32'h8000_0001);
      end
   end
`endif   

   // Gearbox and reset circuitry.
  Clockworks
    // #(.SLOW(21)) // Divide clock frequency by 2^21
  CW(
    .CLK(CLK),
    .RESET(RESET),
    .clk(clk),
    .resetn(resetn)
  );
   

endmodule